package mac_int32p;
typedef struct {Bit#(1) sum;
		Bit#(1) cout;} Adder_output deriving(Bits, Eq); 
typedef struct {Bit#(16) out1;
		Bit#(16) out2;}  Wm_output deriving(Bits, Eq);

import SpecialFIFOs :: *;
import FIFOF :: *;
import DReg :: *;

interface Mac_int_ifc;
	method Action mac_int_input(Bit#(8) inp_1, Bit#(8) inp_2, Bit#(32) inp_3);
	method Bit#(32) mac_int_output();
endinterface : Mac_int_ifc

interface Csa_ifc;
	method Action csa_input(Bit#(32) csa_inp1, Bit#(32) csa_inp2, Bit#(32) csa_inp3);
	method ActionValue#(Bit#(32)) csa_output();
endinterface : Csa_ifc

interface Rca_ifc;
	method Action rca_input(Bit#(32) rca_inp1, Bit#(32) rca_inp2);
	method ActionValue#(Bit#(32)) rca_output();
endinterface : Rca_ifc

interface Wallace_multiplier_ifc;
	method Action wallace_input(Bit#(8) wm_inp1, Bit#(8) wm_inp2);
	method ActionValue#(Bit#(16)) wallace_output();
endinterface : Wallace_multiplier_ifc


module mk_wallace_multiplier(Wallace_multiplier_ifc);

	Csa_ifc csa_unit <- mk_carry_save_adder;
	
	//Partial Product FIFOs
	FIFOF#(Bit#(8)) ff_p00 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p01 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p02 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p03 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p04 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p05 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p06 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_p07 <- mkPipelineFIFOF();
	
	//Level 1 FIFOs
	FIFOF#(Bit#(15)) ff_p10 <- mkPipelineFIFOF();
	FIFOF#(Bit#(13)) ff_p11 <- mkPipelineFIFOF();
	FIFOF#(Bit#(9)) ff_p12 <- mkPipelineFIFOF();
	FIFOF#(Bit#(7)) ff_p13 <- mkPipelineFIFOF();
	FIFOF#(Bit#(3)) ff_p14 <- mkPipelineFIFOF();
	FIFOF#(Bit#(1)) ff_p15 <- mkPipelineFIFOF();
	
	//Level 2 FIFOs
	FIFOF#(Bit#(16)) ff_p20 <- mkPipelineFIFOF();
	FIFOF#(Bit#(12)) ff_p21 <- mkPipelineFIFOF();
	FIFOF#(Bit#(7)) ff_p22 <- mkPipelineFIFOF();
	FIFOF#(Bit#(3)) ff_p23 <- mkPipelineFIFOF();
	
	//Level 3 FIFOs
	FIFOF#(Bit#(16)) ff_p30 <- mkPipelineFIFOF();
	FIFOF#(Bit#(12)) ff_p31 <- mkPipelineFIFOF();
	FIFOF#(Bit#(3)) ff_p32 <- mkPipelineFIFOF();
	
	//Level 4 FIFO
	FIFOF#(Bit#(16)) ff_out <- mkPipelineFIFOF();

	function Adder_output half_adder(Bit#(1) ha_inp1, Bit#(1) ha_inp2);
		Bit#(1) ha_sum  = ha_inp1 ^ ha_inp2;
		Bit#(1) ha_cout = ha_inp1 & ha_inp2;
		Adder_output ha_out = Adder_output{sum: ha_sum, cout: ha_cout};
		return ha_out;
	endfunction : half_adder
	
	function Adder_output full_adder(Bit#(1) f_inp1, Bit#(1) f_inp2, Bit#(1) f_cin);
		Bit#(1) f_sum  = f_inp1 ^ f_inp2 ^ f_cin;
		Bit#(1) f_cout = (f_inp1 & f_inp2) | (f_inp1 & f_cin) | (f_inp2 & f_cin);
		Adder_output f_out = Adder_output{sum: f_sum, cout: f_cout};
		return f_out;
	endfunction : full_adder
	

	rule level_1;
	
		Bit#(8) rg_p00 = ff_p00.first;
		Bit#(8) rg_p01 = ff_p01.first;
		Bit#(8) rg_p02 = ff_p02.first;
		Bit#(8) rg_p03 = ff_p03.first;
		Bit#(8) rg_p04 = ff_p04.first;
		Bit#(8) rg_p05 = ff_p05.first;
		Bit#(8) rg_p06 = ff_p06.first;
		Bit#(8) rg_p07 = ff_p07.first;
	
		Bit#(15) w10 = 0;
		Bit#(13) w11 = 0;
		Bit#(9) w12 = 0;
		Bit#(7) w13 = 0;
		Bit#(3) w14 = 0;
		Bit#(1) w15 = 0;
		
		w10[0] = rg_p00[0];
		let half_adder1 = half_adder(rg_p00[1], rg_p01[0]);
		w10[1] = half_adder1.sum;
		w10[2] = half_adder1.cout;
		let full_adder1 = full_adder(rg_p00[2], rg_p01[1], rg_p02[0]);
		w11[0] = full_adder1.sum;
		w10[3] = full_adder1.cout;
		let full_adder2 = full_adder(rg_p00[3], rg_p01[2], rg_p02[1]);
		w11[1] = full_adder2.sum;
		w10[4] = full_adder2.cout;
		w12[0] = rg_p03[0];
		let full_adder3 = full_adder(rg_p00[4], rg_p01[3], rg_p02[2]);
		w11[2] = full_adder3.sum;
		w10[5] = full_adder3.cout;
		let half_adder2 = half_adder(rg_p03[1], rg_p04[0]);
		w12[1] = half_adder2.sum;
		w11[3] = half_adder2.cout;
		let full_adder4 = full_adder(rg_p00[5], rg_p01[4], rg_p02[3]);
		w12[2] = full_adder4.sum;
		w10[6] = full_adder4.cout;
		let full_adder5 = full_adder(rg_p03[2], rg_p04[1], rg_p05[0]);
		w13[0] = full_adder5.sum;
		w11[4] = full_adder5.cout;
		let full_adder6 = full_adder(rg_p00[6], rg_p01[5], rg_p02[4]);
		w12[3] = full_adder6.sum;
		w10[7] = full_adder6.cout;
		let full_adder7 = full_adder(rg_p03[3], rg_p04[2], rg_p05[1]);
		w13[1] = full_adder7.sum;
		w11[5] = full_adder7.cout;
		w14[0] = rg_p06[0];
		let full_adder8 = full_adder(rg_p00[7], rg_p01[6], rg_p02[5]);
		w12[4] = full_adder8.sum;
		w10[8] = full_adder8.cout;
		let full_adder9 = full_adder(rg_p03[4], rg_p04[3], rg_p05[2]);
		w13[2] = full_adder9.sum;
		w11[6] = full_adder9.cout;
		let half_adder3 = half_adder(rg_p06[1], rg_p07[0]);
		w14[1] = half_adder3.sum;
		w12[5] = half_adder3.cout;		
		let full_adder10 = full_adder(rg_p01[7], rg_p02[6], rg_p03[5]);
		w13[3] = full_adder10.sum;
		w10[9] = full_adder10.cout;
		let full_adder11 = full_adder(rg_p04[4], rg_p05[3], rg_p06[2]);
		w14[2] = full_adder11.sum;
		w11[7] = full_adder11.cout;
		w15    = rg_p07[1];
		let full_adder12 = full_adder(rg_p02[7], rg_p03[6], rg_p04[5]);
		w12[6] = full_adder12.sum;
		w10[10] = full_adder12.cout;
		let full_adder13 = full_adder(rg_p05[4], rg_p06[3], rg_p07[2]);
		w13[4] = full_adder13.sum;
		w11[8] = full_adder13.cout;
		let full_adder14 = full_adder(rg_p03[7], rg_p04[6], rg_p05[5]);
		w12[7] = full_adder14.sum;
		w10[11] = full_adder14.cout;
		let half_adder4 = half_adder(rg_p06[4], rg_p07[3]);
		w13[5] = half_adder4.sum;
		w11[9] = half_adder4.cout;
		let full_adder15 = full_adder(rg_p04[7], rg_p05[6], rg_p06[5]);
		w12[8] = full_adder15.sum;
		w10[12] = full_adder15.cout;
		w13[6] = rg_p07[4];
		let full_adder16 = full_adder(rg_p05[7], rg_p06[6], rg_p07[5]);
		w11[10] = full_adder16.sum;
		w10[13] = full_adder16.cout;
		let half_adder5 = half_adder(rg_p06[7], rg_p07[6]);
		w11[11] = half_adder5.sum;
		w10[14] = half_adder5.cout;
		w11[12] = rg_p07[7];
		
		ff_p10.enq(w10);
		ff_p11.enq(w11);
		ff_p12.enq(w12);
		ff_p13.enq(w13);
		ff_p14.enq(w14);
		ff_p15.enq(w15);
		
		ff_p00.deq;
		ff_p01.deq;
		ff_p02.deq;
		ff_p03.deq;
		ff_p04.deq;
		ff_p05.deq;
		ff_p06.deq;
		ff_p07.deq;

	endrule : level_1		

	rule level_2;
	
		Bit#(15) rg_p10  = ff_p10.first;
		Bit#(13) rg_p11  = ff_p11.first;
		Bit#(9) rg_p12   = ff_p12.first;
		Bit#(7) rg_p13   = ff_p13.first;
		Bit#(3) rg_p14   = ff_p14.first;
		Bit#(1) rg_p15   = ff_p15.first;
	
		Bit#(16) w20 = 0; 
		Bit#(12) w21 = 0; 
		Bit#(7) w22 = 0; 
		Bit#(3) w23 = 0;   
	
		w20[0] = rg_p10[0];
		w20[1] = rg_p10[1];
		let half_adder1 = half_adder(rg_p10[2], rg_p11[0]);
		w20[2] = half_adder1.sum;
		w20[3] = half_adder1.cout;
		let full_adder1 = full_adder(rg_p10[3], rg_p11[1], rg_p12[0]);
		w21[0] = full_adder1.sum;
		w20[4] = full_adder1.cout;
		let full_adder2 = full_adder(rg_p10[4], rg_p11[2], rg_p12[1]);
		w21[1] = full_adder2.sum;
		w20[5] = full_adder2.cout;
		let full_adder3 = full_adder(rg_p10[5], rg_p11[3], rg_p12[2]);
		w21[2] = full_adder3.sum;
		w20[6] = full_adder3.cout;
		w22[0] = rg_p13[0];
		let full_adder4 = full_adder(rg_p10[6], rg_p11[4], rg_p12[3]);
		w21[3] = full_adder4.sum;
		w20[7] = full_adder4.cout;
		let half_adder2 = half_adder(rg_p13[1], rg_p14[0]);
		w22[1] = half_adder2.sum;
		w21[4] = half_adder2.cout;
		let full_adder5 = full_adder(rg_p10[7], rg_p11[5], rg_p12[4]);
		w22[2] = full_adder5.sum;
		w20[8] = full_adder5.cout;
		let half_adder3 = half_adder(rg_p13[2], rg_p14[1]);
		w23[0] = half_adder3.sum;
		w21[5] = half_adder3.cout;
		let full_adder6 = full_adder(rg_p10[8], rg_p11[6], rg_p12[5]);
		w22[3] = full_adder6.sum;
		w20[9] = full_adder6.cout;
		let full_adder7 = full_adder(rg_p13[3], rg_p14[2], rg_p15);
		w23[1] = full_adder7.sum;
		w21[6] = full_adder7.cout;
		let full_adder8 = full_adder(rg_p10[9], rg_p11[7], rg_p12[6]);
		w22[4] = full_adder8.sum;
		w20[10] = full_adder8.cout;
		w23[2] = rg_p13[4];
		let full_adder9 = full_adder(rg_p10[10], rg_p11[8], rg_p12[7]);
		w21[7] = full_adder9.sum;
		w20[11] = full_adder9.cout;
		w22[5] = rg_p13[5];
		let full_adder10 = full_adder(rg_p10[11], rg_p11[9], rg_p12[8]);
		w21[8] = full_adder10.sum;
		w20[12] = full_adder10.cout;
		w22[6] = rg_p13[6];
		let half_adder4 = half_adder(rg_p10[12], rg_p11[10]);
		w21[9] = half_adder4.sum;
		w20[13] = half_adder4.cout;
		let half_adder5 = half_adder(rg_p10[13], rg_p11[11]);
		w21[10] = half_adder5.sum;
		w20[14] = half_adder5.cout;
		let half_adder6 = half_adder(rg_p10[14], rg_p11[12]);
		w21[11] = half_adder6.sum;
		w20[15] = half_adder6.cout;
		
		ff_p20.enq(w20);
		ff_p21.enq(w21);
		ff_p22.enq(w22);
		ff_p23.enq(w23);
		
		ff_p10.deq;
		ff_p11.deq;
		ff_p12.deq;
		ff_p13.deq;
		ff_p14.deq;
		ff_p15.deq;
		
	endrule : level_2

	rule level_3;
	
		Bit#(16) rg_p20  = ff_p20.first;
		Bit#(12) rg_p21  = ff_p21.first;
		Bit#(7) rg_p22   = ff_p22.first;
		Bit#(3) rg_p23   = ff_p23.first;
	
		Bit#(16) w30 = 0;
		Bit#(12) w31 = 0;
		Bit#(3) w32 = 0;

		w30[0] = rg_p20[0];
		w30[1] = rg_p20[1];
		w30[2] = rg_p20[2];
		let half_adder1 = half_adder(rg_p20[3], rg_p21[0]);
		w30[3] = half_adder1.sum;
		w30[4] = half_adder1.cout;		
		let half_adder2 = half_adder(rg_p20[4], rg_p21[1]);
		w31[0] = half_adder2.sum;
		w30[5] = half_adder2.cout;
		let full_adder1 = full_adder(rg_p20[5], rg_p21[2], rg_p22[0]);
		w31[1] = full_adder1.sum;
		w30[6] = full_adder1.cout;
		let full_adder2 = full_adder(rg_p20[6], rg_p21[3], rg_p22[1]);
		w31[2] = full_adder2.sum;
		w30[7] = full_adder2.cout;
		let full_adder3 = full_adder(rg_p20[7], rg_p21[4], rg_p22[2]);
		w31[3] = full_adder3.sum;
		w30[8] = full_adder3.cout;
		w32[0] = rg_p23[0];
		let full_adder4 = full_adder(rg_p20[8], rg_p21[5], rg_p22[3]);
		w31[4] = full_adder4.sum;
		w30[9] = full_adder4.cout;
		w32[1] = rg_p23[1];
		let full_adder5 = full_adder(rg_p20[9], rg_p21[6], rg_p22[4]);
		w31[5] = full_adder5.sum;
		w30[10] = full_adder5.cout;
		w32[2] = rg_p23[2];
		let full_adder6 = full_adder(rg_p20[10], rg_p21[7], rg_p22[5]);
		w31[6] = full_adder6.sum;
		w30[11] = full_adder6.cout;
		let full_adder7 = full_adder(rg_p20[11], rg_p21[8], rg_p22[6]);
		w31[7] = full_adder7.sum;
		w30[12] = full_adder7.cout;
		let half_adder3 = half_adder(rg_p20[12], rg_p21[9]);
		w31[8] = half_adder3.sum;
		w30[13] = half_adder3.cout;
		let half_adder4 = half_adder(rg_p20[13], rg_p21[10]);
		w31[9] = half_adder4.sum;
		w30[14] = half_adder4.cout;
		let half_adder5 = half_adder(rg_p20[14], rg_p21[11]);
		w31[10] = half_adder5.sum;
		w30[15] = half_adder5.cout;
		w31[11] = rg_p20[15];
		
		ff_p30.enq(w30);
		ff_p31.enq(w31);
		ff_p32.enq(w32);		
		
		ff_p20.deq;
		ff_p21.deq;
		ff_p22.deq;
		ff_p23.deq;
	
	endrule : level_3

	rule level_4;
	
		Bit#(16) rg_p30  = ff_p30.first;
		Bit#(12) rg_p31  = ff_p31.first;
		Bit#(3) rg_p32   = ff_p32.first;
	
		Bit#(16) w40 = 0;
		Bit#(16) w41 = 0;
	
		w40[0] = rg_p30[0];
		w40[1] = rg_p30[1];
		w40[2] = rg_p30[2];
		w40[3] = rg_p30[3];
		let half_adder1 = half_adder(rg_p30[4], rg_p31[0]);
		w40[4] = half_adder1.sum;
		w40[5] = half_adder1.cout;		
		let half_adder2 = half_adder(rg_p30[5], rg_p31[1]);
		w41[5] = half_adder2.sum;
		w40[6] = half_adder2.cout;
		let half_adder3 = half_adder(rg_p30[6], rg_p31[2]);
		w41[6] = half_adder3.sum;
		w40[7] = half_adder3.cout;
		let full_adder1 = full_adder(rg_p30[7], rg_p31[3], rg_p32[0]);
		w41[7] = full_adder1.sum;
		w40[8] = full_adder1.cout;
		let full_adder2 = full_adder(rg_p30[8], rg_p31[4], rg_p32[1]);
		w41[8] = full_adder2.sum;
		w40[9] = full_adder2.cout;
		let full_adder3 = full_adder(rg_p30[9], rg_p31[5], rg_p32[2]);
		w41[9] = full_adder3.sum;
		w40[10] = full_adder3.cout;
		let half_adder4 = half_adder(rg_p30[10], rg_p31[6]);
		w41[10] = half_adder4.sum;
		w40[11] = half_adder4.cout;
		let half_adder5 = half_adder(rg_p30[11], rg_p31[7]);
		w41[11] = half_adder5.sum;
		w40[12] = half_adder5.cout;
		let half_adder6 = half_adder(rg_p30[12], rg_p31[8]);
		w41[12] = half_adder6.sum;
		w40[13] = half_adder6.cout;
		let half_adder7 = half_adder(rg_p30[13], rg_p31[9]);
		w41[13] = half_adder7.sum;
		w40[14] = half_adder7.cout;
		let half_adder8 = half_adder(rg_p30[14], rg_p31[10]);
		w41[14] = half_adder8.sum;
		w40[15] = half_adder8.cout;
		let half_adder9 = half_adder(rg_p30[15], rg_p31[11]);
		w41[15] = half_adder9.sum;
		//rg_p41[16] <= half_adder(rg_p30[15], rg_p31[11]).cout;
		
		csa_unit.csa_input(signExtend(w40), signExtend(w41), signExtend(16'b1000000100000000));
		
		
		ff_p30.deq;
		ff_p31.deq;
		ff_p32.deq;		

	endrule : level_4
	
	rule endresult;
	
		Bit#(32) temp <- csa_unit.csa_output();
		Bit#(16) result = truncate(temp);
		ff_out.enq(result);
		
	endrule : endresult

	method Action wallace_input(Bit#(8) wm_inp1, Bit#(8) wm_inp2);
	
		
		Bit#(8) pp0 = (wm_inp1 & {wm_inp2[0], wm_inp2[0], wm_inp2[0], wm_inp2[0], wm_inp2[0], wm_inp2[0], wm_inp2[0], wm_inp2[0]});
		pp0[7] = ~pp0[7];
		Bit#(8) pp1 = (wm_inp1 & {wm_inp2[1], wm_inp2[1], wm_inp2[1], wm_inp2[1], wm_inp2[1], wm_inp2[1], wm_inp2[1], wm_inp2[1]});
		pp1[7] = ~pp1[7];
		Bit#(8) pp2 = (wm_inp1 & {wm_inp2[2], wm_inp2[2], wm_inp2[2], wm_inp2[2], wm_inp2[2], wm_inp2[2], wm_inp2[2], wm_inp2[2]});
		pp2[7] = ~pp2[7];
		Bit#(8) pp3 = (wm_inp1 & {wm_inp2[3], wm_inp2[3], wm_inp2[3], wm_inp2[3], wm_inp2[3], wm_inp2[3], wm_inp2[3], wm_inp2[3]});
		pp3[7] = ~pp3[7];
		Bit#(8) pp4 = (wm_inp1 & {wm_inp2[4], wm_inp2[4], wm_inp2[4], wm_inp2[4], wm_inp2[4], wm_inp2[4], wm_inp2[4], wm_inp2[4]});
		pp4[7] = ~pp4[7];
		Bit#(8) pp5 = (wm_inp1 & {wm_inp2[5], wm_inp2[5], wm_inp2[5], wm_inp2[5], wm_inp2[5], wm_inp2[5], wm_inp2[5], wm_inp2[5]});
		pp5[7] = ~pp5[7];
		Bit#(8) pp6 = (wm_inp1 & {wm_inp2[6], wm_inp2[6], wm_inp2[6], wm_inp2[6], wm_inp2[6], wm_inp2[6], wm_inp2[6], wm_inp2[6]});
		pp6[7] = ~pp6[7];
		Bit#(8) pp7 = (wm_inp1 & {wm_inp2[7], wm_inp2[7], wm_inp2[7], wm_inp2[7], wm_inp2[7], wm_inp2[7], wm_inp2[7], wm_inp2[7]});
		pp7 = ~pp7;
		pp7[7] = ~pp7[7];
		
		ff_p00.enq(pp0);
		ff_p01.enq(pp1);
		ff_p02.enq(pp2);
		ff_p03.enq(pp3);
		ff_p04.enq(pp4);
		ff_p05.enq(pp5);
		ff_p06.enq(pp6);
		ff_p07.enq(pp7);
		
	endmethod : wallace_input
	method ActionValue#(Bit#(16)) wallace_output();
		Bit#(16) result = ff_out.first;
		ff_out.deq;
		return result;
	endmethod : wallace_output
endmodule : mk_wallace_multiplier


module mk_ripple_carry_adder(Rca_ifc);
	
	FIFOF#(Bit#(32)) ff_inp1 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_inp2 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_out <- mkPipelineFIFOF();

	rule addition;
	
		Bit#(32) rg_inp1 = ff_inp1.first;
		Bit#(32) rg_inp2 = ff_inp2.first;
		Bit#(32) sum   = 0;
		Bit#(33) carry = 0;
		for(Integer i = 0; i < 32; i = i + 1)begin
			sum[i] = rg_inp1[i] ^ rg_inp2[i] ^ carry[i];
			carry[i+1] = (rg_inp1[i] & rg_inp2[i]) | (rg_inp1[i] & carry[i]) | (rg_inp2[i] & carry[i]);
		end
		ff_out.enq(sum);
		ff_inp1.deq;
		ff_inp2.deq;
	endrule : addition
	
	method Action rca_input(Bit#(32) rca_inp1, Bit#(32) rca_inp2);
		ff_inp1.enq(rca_inp1);
		ff_inp2.enq(rca_inp2);
	endmethod : rca_input
	method ActionValue#(Bit#(32)) rca_output();
		let rg_out = ff_out.first;
		ff_out.deq;
		return rg_out;
	endmethod : rca_output
endmodule : mk_ripple_carry_adder

module mk_carry_save_adder(Csa_ifc);
		
	Rca_ifc ripple_carry_adder <- mk_ripple_carry_adder;
	
	
	FIFOF#(Bit#(32)) ff_inp1 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_inp2 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_inp3 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_out <- mkPipelineFIFOF();
		
	rule calculation;
	
		Bit#(32) rg_inp1 = ff_inp1.first;
		Bit#(32) rg_inp2 = ff_inp2.first;
		Bit#(32) rg_inp3 = ff_inp3.first;
		
		Bit#(32) sum = 0;
		Bit#(32) carry = 0;
		for(Integer i = 0; i < 32; i = i+1)begin
			sum[i] = (rg_inp1[i] ^ rg_inp2[i] ^ rg_inp3[i]);
			carry[i] = (rg_inp1[i] & rg_inp2[i]) | (rg_inp1[i] & rg_inp3[i]) | (rg_inp2[i] & rg_inp3[i]);
		end
		carry = carry << 1;
		ripple_carry_adder.rca_input(sum, carry);
		ff_inp1.deq;
		ff_inp2.deq;
		ff_inp3.deq;
	endrule : calculation
	rule result;
		Bit#(32) rg_out <- ripple_carry_adder.rca_output();
		ff_out.enq(rg_out);
	endrule : result

	method Action csa_input(Bit#(32) csa_inp1, Bit#(32) csa_inp2, Bit#(32) csa_inp3);
		ff_inp1.enq(csa_inp1);
		ff_inp2.enq(csa_inp2);
		ff_inp3.enq(csa_inp3);
	endmethod : csa_input
	method ActionValue#(Bit#(32)) csa_output();
		let rg_out = ff_out.first;
		ff_out.deq;
		return rg_out;
	endmethod : csa_output

endmodule : mk_carry_save_adder

(*synthesize*)
module mk_mac_int(Mac_int_ifc);

	Wallace_multiplier_ifc wallace_multiplier_unit <- mk_wallace_multiplier;
	Csa_ifc carry_save_adder_unit <- mk_carry_save_adder;

	
	FIFOF#(Bit#(8)) ff_inp_1 <- mkPipelineFIFOF();
	FIFOF#(Bit#(8)) ff_inp_2 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_inp_3 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_inp_3_1 <- mkPipelineFIFOF();
	FIFOF#(Bit#(32)) ff_out <- mkPipelineFIFOF();

	Reg#(Bit#(32)) out <- mkReg(0);
	Reg#(Bool) result_ready <- mkDReg(False);
	
	rule multiplication;
		Bit#(8) rg_inp_1 = ff_inp_1.first;
		Bit#(8) rg_inp_2 = ff_inp_2.first;
		ff_inp_3_1.enq(ff_inp_3.first);
		wallace_multiplier_unit.wallace_input(rg_inp_1, rg_inp_2);
		ff_inp_1.deq;
		ff_inp_2.deq;
		ff_inp_3.deq;
	endrule : multiplication

	rule accumulation;
		Bit#(16) multiplication_ouput <-  wallace_multiplier_unit.wallace_output();
		Bit#(32) input_1 = signExtend(multiplication_ouput);
		Bit#(32) rg_inp_3 = ff_inp_3_1.first;
		carry_save_adder_unit.csa_input(input_1, 32'b0, rg_inp_3);
		ff_inp_3_1.deq;
	endrule : accumulation 

	rule result;
		Bit#(32) rg_out <- carry_save_adder_unit.csa_output();
		out <= rg_out;
		result_ready <= True;
	endrule : result
	
	method Action mac_int_input(Bit#(8) inp_1, Bit#(8) inp_2, Bit#(32) inp_3);
		ff_inp_1.enq(inp_1);
		ff_inp_2.enq(inp_2);
		ff_inp_3.enq(inp_3);
	endmethod : mac_int_input

	method Bit#(32) mac_int_output() if(result_ready);
		Bit#(32) rg_out = out;
		return rg_out;
	endmethod : mac_int_output
endmodule : mk_mac_int
endpackage : mac_int32p


